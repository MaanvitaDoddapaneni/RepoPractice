-- library declaration
-- entity
-- architecture
